
module hps_reset (
	source,
	source_clk);	

	output	[2:0]	source;
	input		source_clk;
endmodule
